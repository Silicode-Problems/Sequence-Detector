//sequence detector for 1011, overlapping

module seq_dec(input wire clk,
                input wire reset,
                input wire in_vl,
                output wire out);
    
   //your code here

endmodule

